import CacheTypes::*;
import Fifo::*;

// TODO: implement message FIFO

module mkMessageFifo(MessageFifo#(n));

endmodule

