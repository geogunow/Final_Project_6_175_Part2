import CacheTypes::*;
import Vector::*;
import MemTypes::*;
import Types::*;
import ProcTypes::*;
import Fifo::*;
import Ehr::*;

// TODO: copy ICache.bsv from project part 1 to here

module mkICache(WideMem mem, ICache ifc);

endmodule

